library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 4;
          addrWidth: natural := 9
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
		  
		  
  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI  : std_logic_vector(3 downto 0) := "0100";
  constant STA  : std_logic_vector(3 downto 0) := "0101";
  constant JMP  : std_logic_vector(3 downto 0) := "0110";
  constant JEQ  : std_logic_vector(3 downto 0) := "0111";
  constant CEQ  : std_logic_vector(3 downto 0) := "1000";
  constant JSR  : std_logic_vector(3 downto 0) := "1001";
  constant RET  : std_logic_vector(3 downto 0) := "1010";

		  
		  
  begin
      -- Palavra de Controle = SelMUX, Habilita_A, Reset_A, Operacao_ULA
      -- Inicializa os endereços:
tmp(0) := "0000000000000";	-- Reset:
tmp(1) := "0101111111110";	-- STA @510
tmp(2) := "0101111111111";	-- STA @511
tmp(3) := "0101111111101";	-- STA @509
tmp(4) := "0100000000000";	-- LDI $0
tmp(5) := "0101000000000";	-- STA @0
tmp(6) := "0101100000010";	-- STA @258
tmp(7) := "0101100000001";	-- STA @257
tmp(8) := "0101100000000";	-- STA @256
tmp(9) := "0101100100000";	-- STA @288
tmp(10) := "0101100100001";	-- STA @289
tmp(11) := "0101100100010";	-- STA @290
tmp(12) := "0101100100011";	-- STA @291
tmp(13) := "0101100100100";	-- STA @292
tmp(14) := "0101100100101";	-- STA @293
tmp(15) := "0101000111111";	-- STA @63
tmp(16) := "0101000111110";	-- STA @62
tmp(17) := "0101000111101";	-- STA @61
tmp(18) := "0101000111100";	-- STA @60
tmp(19) := "0101000111011";	-- STA @59
tmp(20) := "0101000111010";	-- STA @58
tmp(21) := "0101000000010";	-- STA @2
tmp(22) := "0101000000011";	-- STA @3
tmp(23) := "0101000000100";	-- STA @4
tmp(24) := "0101000000101";	-- STA @5
tmp(25) := "0101000000110";	-- STA @6
tmp(26) := "0101000000111";	-- STA @7
tmp(27) := "0100000000001";	-- LDI $1
tmp(28) := "0101000000001";	-- STA @1
tmp(29) := "0100000001010";	-- LDI $10
tmp(30) := "0101000001010";	-- STA @10
tmp(31) := "0000000000000";	-- Inicio:
tmp(32) := "0001101100001";	-- LDA @353
tmp(33) := "1000000000000";	-- CEQ @0
tmp(34) := "0111000011111";	-- JEQ @Inicio
tmp(35) := "1001001000010";	-- JSR @Limite
tmp(36) := "0001000000000";	-- LDA @0
tmp(37) := "0101100100000";	-- STA @288
tmp(38) := "0101100100001";	-- STA @289
tmp(39) := "0101100100010";	-- STA @290
tmp(40) := "0101100100011";	-- STA @291
tmp(41) := "0101100100100";	-- STA @292
tmp(42) := "0101100100101";	-- STA @293
tmp(43) := "0101111111110";	-- STA @510
tmp(44) := "0000000000000";	-- Contador:
tmp(45) := "0000000000000";	-- NOP
tmp(46) := "0001101100000";	-- LDA @352
tmp(47) := "1000000000000";	-- CEQ @0
tmp(48) := "0111001000000";	-- JEQ @LOOP
tmp(49) := "1001001111011";	-- JSR @Incrementa
tmp(50) := "0000000000000";	-- NOP
tmp(51) := "0001000000010";	-- LDA @2
tmp(52) := "0101100100000";	-- STA @288
tmp(53) := "0001000000011";	-- LDA @3
tmp(54) := "0101100100001";	-- STA @289
tmp(55) := "0001000000100";	-- LDA @4
tmp(56) := "0101100100010";	-- STA @290
tmp(57) := "0001000000101";	-- LDA @5
tmp(58) := "0101100100011";	-- STA @291
tmp(59) := "0001000000110";	-- LDA @6
tmp(60) := "0101100100100";	-- STA @292
tmp(61) := "0001000000111";	-- LDA @7
tmp(62) := "0101100100101";	-- STA @293
tmp(63) := "1001010110100";	-- JSR @Comparador
tmp(64) := "0000000000000";	-- LOOP:
tmp(65) := "0110000101100";	-- JMP @Contador
tmp(66) := "0000000000000";	-- Limite:
tmp(67) := "0101111111110";	-- STA @510
tmp(68) := "0000000000000";	-- Unidade:
tmp(69) := "0001101000000";	-- LDA @320
tmp(70) := "0101100100000";	-- STA @288
tmp(71) := "0001101100001";	-- LDA @353
tmp(72) := "1000000000000";	-- CEQ @0
tmp(73) := "0111001000100";	-- JEQ @Unidade
tmp(74) := "0101111111110";	-- STA @510
tmp(75) := "0001101000000";	-- LDA @320
tmp(76) := "0101000111111";	-- STA @63
tmp(77) := "0000000000000";	-- Dezena:
tmp(78) := "0001101000000";	-- LDA @320
tmp(79) := "0101100100001";	-- STA @289
tmp(80) := "0001101100001";	-- LDA @353
tmp(81) := "1000000000000";	-- CEQ @0
tmp(82) := "0111001001101";	-- JEQ @Dezena
tmp(83) := "0101111111110";	-- STA @510
tmp(84) := "0001101000000";	-- LDA @320
tmp(85) := "0101000111110";	-- STA @62
tmp(86) := "0000000000000";	-- Centena:
tmp(87) := "0001101000000";	-- LDA @320
tmp(88) := "0101100100010";	-- STA @290
tmp(89) := "0001101100001";	-- LDA @353
tmp(90) := "1000000000000";	-- CEQ @0
tmp(91) := "0111001010110";	-- JEQ @Centena
tmp(92) := "0101111111110";	-- STA @510
tmp(93) := "0001101000000";	-- LDA @320
tmp(94) := "0101000111101";	-- STA @61
tmp(95) := "0000000000000";	-- Milhar:
tmp(96) := "0001101000000";	-- LDA @320
tmp(97) := "0101100100011";	-- STA @291
tmp(98) := "0001101100001";	-- LDA @353
tmp(99) := "1000000000000";	-- CEQ @0
tmp(100) := "0111001011111";	-- JEQ @Milhar
tmp(101) := "0101111111110";	-- STA @510
tmp(102) := "0001101000000";	-- LDA @320
tmp(103) := "0101000111100";	-- STA @60
tmp(104) := "0000000000000";	-- DezMilhar:
tmp(105) := "0001101000000";	-- LDA @320
tmp(106) := "0101100100100";	-- STA @292
tmp(107) := "0001101100001";	-- LDA @353
tmp(108) := "1000000000000";	-- CEQ @0
tmp(109) := "0111001101000";	-- JEQ @DezMilhar
tmp(110) := "0101111111110";	-- STA @510
tmp(111) := "0001101000000";	-- LDA @320
tmp(112) := "0101000111011";	-- STA @59
tmp(113) := "0000000000000";	-- CenMilhar:
tmp(114) := "0001101000000";	-- LDA @320
tmp(115) := "0101100100101";	-- STA @293
tmp(116) := "0001101100001";	-- LDA @353
tmp(117) := "1000000000000";	-- CEQ @0
tmp(118) := "0111001110001";	-- JEQ @CenMilhar
tmp(119) := "0101111111110";	-- STA @510
tmp(120) := "0001101000000";	-- LDA @320
tmp(121) := "0101000111010";	-- STA @58
tmp(122) := "1010000000000";	-- RET
tmp(123) := "0000000000000";	-- Incrementa:
tmp(124) := "0101111111111";	-- STA @511
tmp(125) := "0001000000010";	-- LDA @2
tmp(126) := "0010000000001";	-- SOMA @1
tmp(127) := "1000000001010";	-- CEQ @10
tmp(128) := "0111010000011";	-- JEQ @Dez
tmp(129) := "0101000000010";	-- STA @2
tmp(130) := "1010000000000";	-- RET
tmp(131) := "0000000000000";	-- Dez:
tmp(132) := "0001000000000";	-- LDA @0
tmp(133) := "0101000000010";	-- STA @2
tmp(134) := "0001000000011";	-- LDA @3
tmp(135) := "0010000000001";	-- SOMA @1
tmp(136) := "1000000001010";	-- CEQ @10
tmp(137) := "0111010001100";	-- JEQ @Cen
tmp(138) := "0101000000011";	-- STA @3
tmp(139) := "1010000000000";	-- RET
tmp(140) := "0000000000000";	-- Cen:
tmp(141) := "0001000000000";	-- LDA @0
tmp(142) := "0101000000011";	-- STA @3
tmp(143) := "0001000000100";	-- LDA @4
tmp(144) := "0010000000001";	-- SOMA @1
tmp(145) := "1000000001010";	-- CEQ @10
tmp(146) := "0111010010101";	-- JEQ @Mil
tmp(147) := "0101000000100";	-- STA @4
tmp(148) := "1010000000000";	-- RET
tmp(149) := "0000000000000";	-- Mil:
tmp(150) := "0001000000000";	-- LDA @0
tmp(151) := "0101000000100";	-- STA @4
tmp(152) := "0001000000101";	-- LDA @5
tmp(153) := "0010000000001";	-- SOMA @1
tmp(154) := "1000000001010";	-- CEQ @10
tmp(155) := "0111010011110";	-- JEQ @DezM
tmp(156) := "0101000000101";	-- STA @5
tmp(157) := "1010000000000";	-- RET
tmp(158) := "0000000000000";	-- DezM:
tmp(159) := "0001000000000";	-- LDA @0
tmp(160) := "0101000000101";	-- STA @5
tmp(161) := "0001000000110";	-- LDA @6
tmp(162) := "0010000000001";	-- SOMA @1
tmp(163) := "1000000001010";	-- CEQ @10
tmp(164) := "0111010100111";	-- JEQ @CenM
tmp(165) := "0101000000110";	-- STA @6
tmp(166) := "1010000000000";	-- RET
tmp(167) := "0000000000000";	-- CenM:
tmp(168) := "0001000000000";	-- LDA @0
tmp(169) := "0101000000110";	-- STA @6
tmp(170) := "0001000000111";	-- LDA @7
tmp(171) := "0010000000001";	-- SOMA @1
tmp(172) := "1000000001010";	-- CEQ @10
tmp(173) := "0111010110000";	-- JEQ @Fim
tmp(174) := "0101000000111";	-- STA @7
tmp(175) := "1010000000000";	-- RET
tmp(176) := "0000000000000";	-- Fim:
tmp(177) := "0001000000000";	-- LDA @0
tmp(178) := "0101000000111";	-- STA @7
tmp(179) := "1010000000000";	-- RET
tmp(180) := "0000000000000";	-- Comparador:
tmp(181) := "0001000111111";	-- LDA @63
tmp(182) := "1000000000010";	-- CEQ @2
tmp(183) := "0111010111001";	-- JEQ @CompDez
tmp(184) := "1010000000000";	-- RET
tmp(185) := "0000000000000";	-- CompDez:
tmp(186) := "0001000111110";	-- LDA @62
tmp(187) := "1000000000011";	-- CEQ @3
tmp(188) := "0111010111110";	-- JEQ @CompCen
tmp(189) := "1010000000000";	-- RET
tmp(190) := "0000000000000";	-- CompCen:
tmp(191) := "0001000111101";	-- LDA @61
tmp(192) := "1000000000100";	-- CEQ @4
tmp(193) := "0111011000011";	-- JEQ @CompMil
tmp(194) := "1010000000000";	-- RET
tmp(195) := "0000000000000";	-- CompMil:
tmp(196) := "0001000111100";	-- LDA @60
tmp(197) := "1000000000101";	-- CEQ @5
tmp(198) := "0111011001000";	-- JEQ @CompDezM
tmp(199) := "1010000000000";	-- RET
tmp(200) := "0000000000000";	-- CompDezM:
tmp(201) := "0001000111011";	-- LDA @59
tmp(202) := "1000000000110";	-- CEQ @6
tmp(203) := "0111011001101";	-- JEQ @CompCenM
tmp(204) := "1010000000000";	-- RET
tmp(205) := "0000000000000";	-- CompCenM:
tmp(206) := "0001000111010";	-- LDA @58
tmp(207) := "1000000000111";	-- CEQ @7
tmp(208) := "0111011010010";	-- JEQ @Acabou
tmp(209) := "1010000000000";	-- RET
tmp(210) := "0000000000000";	-- Acabou:
tmp(211) := "0100000000001";	-- LDI @1
tmp(212) := "0101100000010";	-- STA @258
tmp(213) := "0101100000001";	-- STA @257
tmp(214) := "0100011111111";	-- LDI $255
tmp(215) := "0101100000000";	-- STA @256
tmp(216) := "0001101100100";	-- LDA @356
tmp(217) := "1000000000000";	-- CEQ @0
tmp(218) := "0111011010010";	-- JEQ @Acabou
tmp(219) := "0110000000000";	-- JMP @Reset





        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;
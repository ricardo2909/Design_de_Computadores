library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 4;
          addrWidth: natural := 9
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
		  
		  
  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI  : std_logic_vector(3 downto 0) := "0100";
  constant STA  : std_logic_vector(3 downto 0) := "0101";
  constant JMP  : std_logic_vector(3 downto 0) := "0110";
  constant JEQ  : std_logic_vector(3 downto 0) := "0111";
  constant CEQ  : std_logic_vector(3 downto 0) := "1000";
  constant JSR  : std_logic_vector(3 downto 0) := "1001";
  constant RET  : std_logic_vector(3 downto 0) := "1010";

		  
		  
  begin
      -- Palavra de Controle = SelMUX, Habilita_A, Reset_A, Operacao_ULA
      -- Inicializa os endereços:
tmp(0) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(1) := x"5" & "00" & '1' & x"FE";	-- STA @510                    	#Limpa leitura KEY1
tmp(2) := x"5" & "00" & '1' & x"FF";	-- STA @511                    	#Limpa leitura KEY0
tmp(3) := x"5" & "00" & '1' & x"FD";	-- STA @509                    	#Limpa leitura Reset    
tmp(4) := x"4" & "00" & '0' & x"01";	-- LDI $1                      	#Carrega 1 no acumulador
tmp(5) := x"5" & "00" & '0' & x"3F";	-- STA @63                     	#Salva 1 no endereço 63 da RAM
tmp(6) := x"4" & "00" & '0' & x"09";	-- LDI $9                      	#Carrega 9 no acumulador
tmp(7) := x"5" & "00" & '0' & x"13";	-- STA @19                     	#Salva 9 no endereço 19 da RAM
tmp(8) := x"4" & "00" & '0' & x"0A";	-- LDI $10                     	#Carrega 10 no acumulador
tmp(9) := x"5" & "00" & '0' & x"14";	-- STA @20                     	#Salva 10 no endereço 20 da RAM
tmp(10) := x"4" & "00" & '0' & x"0B";	-- LDI $11                     	#Carrega 11 no acumulador
tmp(11) := x"5" & "00" & '0' & x"15";	-- STA @21                     	#Salva 11 no endereço 21 da RAM
tmp(12) := x"4" & "00" & '0' & x"0C";	-- LDI $12                     	#Carrega 12 no acumulador
tmp(13) := x"5" & "00" & '0' & x"16";	-- STA @22                     	#Salva 12 no endereço 22 da RAM
tmp(14) := x"4" & "00" & '0' & x"0D";	-- LDI $13                     	#Carrega 13 no acumulador
tmp(15) := x"5" & "00" & '0' & x"17";	-- STA @23                     	#Salva 13 no endereço 23 da RAM
tmp(16) := x"4" & "00" & '0' & x"0E";	-- LDI $14                     	#Carrega 14 no acumulador
tmp(17) := x"5" & "00" & '0' & x"18";	-- STA @24                     	#Salva 14 no endereço 24 da RAM
tmp(18) := x"4" & "00" & '0' & x"0F";	-- LDI $15                     	#Carrega 15 no acumulador
tmp(19) := x"5" & "00" & '0' & x"19";	-- STA @25                     	#Salva 15 no endereço 25 da RAM
tmp(20) := x"4" & "00" & '0' & x"00";	-- LDI $0                      	#Carrega 0 no acumulador
tmp(21) := x"5" & "00" & '0' & x"3E";	-- STA @62                     	#Salva 0 no endereço 62 da RAM
tmp(22) := x"5" & "00" & '1' & x"02";	-- STA @258                    	#Apaga o LED 9
tmp(23) := x"5" & "00" & '1' & x"01";	-- STA @257                    	#Apaga o LED 8
tmp(24) := x"5" & "00" & '1' & x"00";	-- STA @256                    	#Apaga o LED 7 a 0 
tmp(25) := x"5" & "00" & '1' & x"20";	-- STA @288                    	#Zera o HEX 0
tmp(26) := x"5" & "00" & '1' & x"21";	-- STA @289                    	#Zera o HEX 1
tmp(27) := x"5" & "00" & '1' & x"22";	-- STA @290                    	#Zera o HEX 2
tmp(28) := x"5" & "00" & '1' & x"23";	-- STA @291                    	#Zera o HEX 3
tmp(29) := x"5" & "00" & '1' & x"24";	-- STA @292                    	#Zera o HEX 4
tmp(30) := x"5" & "00" & '1' & x"25";	-- STA @293                    	#Zera o HEX 5
tmp(31) := x"5" & "00" & '0' & x"00";	-- STA @0                      	#Zera o endereço 0 da RAM (Limite das unidades)
tmp(32) := x"5" & "00" & '0' & x"01";	-- STA @1                      	#Zera o endereço 1 da RAM (Limite das dezenas)
tmp(33) := x"5" & "00" & '0' & x"02";	-- STA @2                      	#Zera o endereço 2 da RAM (Limite das centenas) 
tmp(34) := x"5" & "00" & '0' & x"03";	-- STA @3                      	#Zera o endereço 3 da RAM (Limite dos milhares) 
tmp(35) := x"5" & "00" & '0' & x"04";	-- STA @4                      	#Zera o endereço 4 da RAM (Limite das dezenas de milhares)
tmp(36) := x"5" & "00" & '0' & x"05";	-- STA @5                      	#Zera o endereço 5 da RAM (Limite das centenas de milhares) 
tmp(37) := x"5" & "00" & '0' & x"0A";	-- STA @10                     	#Zera o endereço 10 da RAM (Valor atual das unidades) 
tmp(38) := x"5" & "00" & '0' & x"0B";	-- STA @11                     	#Zera o endereço 11 da RAM (Valor atual das dezenas)
tmp(39) := x"5" & "00" & '0' & x"0C";	-- STA @12                     	#Zera o endereço 12 da RAM (Valor atual das centenas)
tmp(40) := x"5" & "00" & '0' & x"0D";	-- STA @13                     	#Zera o endereço 13 da RAM (Valor atual dos milhares)
tmp(41) := x"5" & "00" & '0' & x"0E";	-- STA @14                     	#Zera o endereço 14 da RAM (Valor atual das dezenas de milhares)
tmp(42) := x"5" & "00" & '0' & x"0F";	-- STA @15                     	#Zera o endereço 15 da RAM (Valor atual das centenas de milhares)
tmp(43) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(44) := x"1" & "00" & '1' & x"61";	-- LDA @353                    	#Carrega o valor do KEY1 no acumulador
tmp(45) := x"8" & "00" & '0' & x"3F";	-- CEQ @63                     	#Compara o valor do KEY1 com 63 (1)
tmp(46) := x"7" & "00" & '0' & x"36";	-- JEQ @54           	#Se o valor do KEY1 for 1, vai para o label SetLim (Setar Limite)
tmp(47) := x"1" & "00" & '1' & x"60";	-- LDA @352                    	#Carrega o valor do KEY0 no acumulador
tmp(48) := x"8" & "00" & '0' & x"3F";	-- CEQ @63                     	#Compara o valor do KEY0 com 63 (1)
tmp(49) := x"7" & "00" & '0' & x"ED";	-- JEQ @237           	#Se o valor do KEY0 for 1, vai para o label Incremento (Incrementar)
tmp(50) := x"1" & "00" & '1' & x"64";	-- LDA @356                    	#Carrega o valor do Reset no acumulador
tmp(51) := x"8" & "00" & '0' & x"3F";	-- CEQ @63                     	#Compara o valor do Reset com 63 (1)
tmp(52) := x"7" & "00" & '0' & x"00";	-- JEQ @0           	#Se o valor do Reset for 1, vai para o label Reset (Reseta o programa)
tmp(53) := x"6" & "00" & '0' & x"2B";	-- JMP @43           	#Se nenhum dos botoes forem clicados, vai para o label Start (Laco principal)
tmp(54) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(55) := x"5" & "00" & '1' & x"FE";	-- STA @510                    	#Limpa leitura KEY1
tmp(56) := x"1" & "00" & '0' & x"00";	-- LDA @0                      	#Carrega o valor do endereço 0 da RAM no acumulador (Limite das unidades)
tmp(57) := x"5" & "00" & '1' & x"20";	-- STA @288                    	#Mostra o valor do acumulador HEX 0 (unidades)
tmp(58) := x"1" & "00" & '0' & x"01";	-- LDA @1                      	#Carrega o valor do endereço 1 da RAM no acumulador (Limite das dezenas)
tmp(59) := x"5" & "00" & '1' & x"21";	-- STA @289                    	#Mostra o valor do acumulador HEX 1 (dezenas)
tmp(60) := x"1" & "00" & '0' & x"02";	-- LDA @2                      	#Carrega o valor do endereço 2 da RAM no acumulador (Limite das centenas)
tmp(61) := x"5" & "00" & '1' & x"22";	-- STA @290                    	#Mostra o valor do acumulador HEX 2 (centenas)
tmp(62) := x"1" & "00" & '0' & x"03";	-- LDA @3                      	#Carrega o valor do endereço 3 da RAM no acumulador (Limite dos milhares)
tmp(63) := x"5" & "00" & '1' & x"23";	-- STA @291                    	#Mostra o valor do acumulador HEX 3 (milhares)
tmp(64) := x"1" & "00" & '0' & x"04";	-- LDA @4                      	#Carrega o valor do endereço 4 da RAM no acumulador (Limite das dezenas de milhares)
tmp(65) := x"5" & "00" & '1' & x"24";	-- STA @292                    	#Mostra o valor do acumulador HEX 4 (dezenas de milhares)
tmp(66) := x"1" & "00" & '0' & x"05";	-- LDA @5                      	#Carrega o valor do endereço 5 da RAM no acumulador (Limite das centenas de milhares)
tmp(67) := x"5" & "00" & '1' & x"25";	-- STA @293                    	#Mostra o valor do acumulador HEX 5 (centenas de milhares)
tmp(68) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(69) := x"1" & "00" & '1' & x"40";	-- LDA @320                    	#Carrega valor das chaves SW0 a SW7 no acumulador
tmp(70) := x"8" & "00" & '0' & x"14";	-- CEQ @20                     	#Compara o valor das chaves SW0 a SW7 com 20 (10)
tmp(71) := x"7" & "00" & '0' & x"55";	-- JEQ @85           	#Se o valor das chaves SW0 a SW7 for 10, vai para o label maxUni (Limite maximo das unidades)
tmp(72) := x"8" & "00" & '0' & x"15";	-- CEQ @21                     	#Compara o valor das chaves SW0 a SW7 com 21 (11)
tmp(73) := x"7" & "00" & '0' & x"55";	-- JEQ @85           	#Se o valor das chaves SW0 a SW7 for 11, vai para o label maxUni (Limite maximo das unidades)
tmp(74) := x"8" & "00" & '0' & x"16";	-- CEQ @22                     	#Compara o valor das chaves SW0 a SW7 com 22 (12)
tmp(75) := x"7" & "00" & '0' & x"55";	-- JEQ @85           	#Se o valor das chaves SW0 a SW7 for 12, vai para o label maxUni (Limite maximo das unidades)
tmp(76) := x"8" & "00" & '0' & x"17";	-- CEQ @23                     	#Compara o valor das chaves SW0 a SW7 com 23 (13)
tmp(77) := x"7" & "00" & '0' & x"55";	-- JEQ @85           	#Se o valor das chaves SW0 a SW7 for 13, vai para o label maxUni (Limite maximo das unidades)
tmp(78) := x"8" & "00" & '0' & x"18";	-- CEQ @24                     	#Compara o valor das chaves SW0 a SW7 com 24 (14)
tmp(79) := x"7" & "00" & '0' & x"55";	-- JEQ @85           	#Se o valor das chaves SW0 a SW7 for 14, vai para o label maxUni (Limite maximo das unidades)
tmp(80) := x"8" & "00" & '0' & x"19";	-- CEQ @25                     	#Compara o valor das chaves SW0 a SW7 com 25 (15)
tmp(81) := x"7" & "00" & '0' & x"55";	-- JEQ @85           	#Se o valor das chaves SW0 a SW7 for 15, vai para o label maxUni (Limite maximo das unidades)
tmp(82) := x"5" & "00" & '1' & x"20";	-- STA @288                    	#Mostra o valor do acumulador HEX 0 (unidades)
tmp(83) := x"5" & "00" & '0' & x"00";	-- STA @0                      	#Salva o valor do acumulador no endereço 0 da RAM (Limite das unidades)
tmp(84) := x"6" & "00" & '0' & x"59";	-- JMP @89           	#Vai para o label UNIOK (Unidades menor que o limite)
tmp(85) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(86) := x"1" & "00" & '0' & x"13";	-- LDA @19                     	#Carrega o endereco 19 da RAM no acumulador (9)
tmp(87) := x"5" & "00" & '1' & x"20";	-- STA @288                    	#Mostra o valor do acumulador HEX 0 (unidades)
tmp(88) := x"5" & "00" & '0' & x"00";	-- STA @0                      	#Salva 9 no endereço 0 da RAM (Limite das unidades)
tmp(89) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(90) := x"1" & "00" & '1' & x"61";	-- LDA @353                    	#Carrega o valor do KEY1 no acumulador
tmp(91) := x"8" & "00" & '0' & x"3E";	-- CEQ @62                     	#Compara o valor do KEY1 com 62 (0)
tmp(92) := x"7" & "00" & '0' & x"44";	-- JEQ @68           	#Se o valor do KEY1 for 0 (nao setou o limite das unidades), vai para o label LimUni (Limite das unidades)
tmp(93) := x"5" & "00" & '1' & x"FE";	-- STA @510                    	#Limpa leitura KEY1
tmp(94) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(95) := x"1" & "00" & '1' & x"40";	-- LDA @320                    	#Carrega valor das chaves SW0 a SW7 no acumulador
tmp(96) := x"8" & "00" & '0' & x"14";	-- CEQ @20                     	#Compara o valor das chaves SW0 a SW7 com 20 (10)
tmp(97) := x"7" & "00" & '0' & x"6F";	-- JEQ @111           	#Se o valor das chaves SW0 a SW7 for 10, vai para o label maxDez (Limite maximo das dezenas)
tmp(98) := x"8" & "00" & '0' & x"15";	-- CEQ @21                     	#Compara o valor das chaves SW0 a SW7 com 21 (11)
tmp(99) := x"7" & "00" & '0' & x"6F";	-- JEQ @111           	#Se o valor das chaves SW0 a SW7 for 11, vai para o label maxDez (Limite maximo das dezenas)
tmp(100) := x"8" & "00" & '0' & x"16";	-- CEQ @22                     	#Compara o valor das chaves SW0 a SW7 com 22 (12)
tmp(101) := x"7" & "00" & '0' & x"6F";	-- JEQ @111           	#Se o valor das chaves SW0 a SW7 for 12, vai para o label maxDez (Limite maximo das dezenas)
tmp(102) := x"8" & "00" & '0' & x"17";	-- CEQ @23                     	#Compara o valor das chaves SW0 a SW7 com 23 (13)
tmp(103) := x"7" & "00" & '0' & x"6F";	-- JEQ @111           	#Se o valor das chaves SW0 a SW7 for 13, vai para o label maxDez (Limite maximo das dezenas)
tmp(104) := x"8" & "00" & '0' & x"18";	-- CEQ @24                     	#Compara o valor das chaves SW0 a SW7 com 24 (14)
tmp(105) := x"7" & "00" & '0' & x"6F";	-- JEQ @111           	#Se o valor das chaves SW0 a SW7 for 14, vai para o label maxDez (Limite maximo das dezenas)
tmp(106) := x"8" & "00" & '0' & x"19";	-- CEQ @25                     	#Compara o valor das chaves SW0 a SW7 com 25 (15)
tmp(107) := x"7" & "00" & '0' & x"6F";	-- JEQ @111           	#Se o valor das chaves SW0 a SW7 for 15, vai para o label maxDez (Limite maximo das dezenas)
tmp(108) := x"5" & "00" & '1' & x"21";	-- STA @289                    	#Mostra o valor do acumulador HEX 1 (dezenas)
tmp(109) := x"5" & "00" & '0' & x"01";	-- STA @1                      	#Salva o valor do acumulador no endereço 1 da RAM (Limite das dezenas)
tmp(110) := x"6" & "00" & '0' & x"73";	-- JMP @115           	#Vai para o label DEZOK (Dezenas menor que o limite)
tmp(111) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(112) := x"1" & "00" & '0' & x"13";	-- LDA @19                     	#Carrega 19 no acumulador
tmp(113) := x"5" & "00" & '1' & x"21";	-- STA @289                    	#Mostra o valor do acumulador HEX 1 (dezenas)
tmp(114) := x"5" & "00" & '0' & x"01";	-- STA @1                      	#Salva 9 no endereço 1 da RAM (Limite das dezenas)
tmp(115) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(116) := x"1" & "00" & '1' & x"61";	-- LDA @353                    	#Carrega o valor do KEY1 no acumulador
tmp(117) := x"8" & "00" & '0' & x"3E";	-- CEQ @62                     	#Compara o valor do KEY1 com 62 (0)
tmp(118) := x"7" & "00" & '0' & x"5E";	-- JEQ @94           	#Se o valor do KEY1 for 0 (nao setou o limite das dezenas), vai para o label LimDez (Limite das dezenas)
tmp(119) := x"5" & "00" & '1' & x"FE";	-- STA @510                    	#Limpa leitura KEY1
tmp(120) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(121) := x"1" & "00" & '1' & x"40";	-- LDA @320                    	#Carrega valor das chaves SW0 a SW7 no acumulador
tmp(122) := x"8" & "00" & '0' & x"14";	-- CEQ @20                     	#Compara o valor das chaves SW0 a SW7 com 20 (10)
tmp(123) := x"7" & "00" & '0' & x"89";	-- JEQ @137           	#Se o valor das chaves SW0 a SW7 for 10, vai para o label maxCen (Limite maximo das centenas)
tmp(124) := x"8" & "00" & '0' & x"15";	-- CEQ @21                     	#Compara o valor das chaves SW0 a SW7 com 21 (11)
tmp(125) := x"7" & "00" & '0' & x"89";	-- JEQ @137           	#Se o valor das chaves SW0 a SW7 for 11, vai para o label maxCen (Limite maximo das centenas)
tmp(126) := x"8" & "00" & '0' & x"16";	-- CEQ @22                     	#Compara o valor das chaves SW0 a SW7 com 22 (12)
tmp(127) := x"7" & "00" & '0' & x"89";	-- JEQ @137           	#Se o valor das chaves SW0 a SW7 for 12, vai para o label maxCen (Limite maximo das centenas)
tmp(128) := x"8" & "00" & '0' & x"17";	-- CEQ @23                     	#Compara o valor das chaves SW0 a SW7 com 23 (13)
tmp(129) := x"7" & "00" & '0' & x"89";	-- JEQ @137           	#Se o valor das chaves SW0 a SW7 for 13, vai para o label maxCen (Limite maximo das centenas)
tmp(130) := x"8" & "00" & '0' & x"18";	-- CEQ @24                     	#Compara o valor das chaves SW0 a SW7 com 24 (14)
tmp(131) := x"7" & "00" & '0' & x"89";	-- JEQ @137           	#Se o valor das chaves SW0 a SW7 for 14, vai para o label maxCen (Limite maximo das centenas)
tmp(132) := x"8" & "00" & '0' & x"19";	-- CEQ @25                     	#Compara o valor das chaves SW0 a SW7 com 25 (15)
tmp(133) := x"7" & "00" & '0' & x"89";	-- JEQ @137           	#Se o valor das chaves SW0 a SW7 for 15, vai para o label maxCen (Limite maximo das centenas)
tmp(134) := x"5" & "00" & '1' & x"22";	-- STA @290                    	#Mostra o valor do acumulador HEX 2 (centenas)
tmp(135) := x"5" & "00" & '0' & x"02";	-- STA @2                      	#Salva o valor do acumulador no endereço 2 da RAM (Limite das centenas)
tmp(136) := x"6" & "00" & '0' & x"8D";	-- JMP @141           	#Vai para o label CENOK (Centenas menor que o limite)
tmp(137) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(138) := x"1" & "00" & '0' & x"13";	-- LDA @19                     	#Carrega 19 no acumulador
tmp(139) := x"5" & "00" & '1' & x"22";	-- STA @290                    	#Mostra o valor do acumulador HEX 2 (centenas)
tmp(140) := x"5" & "00" & '0' & x"02";	-- STA @2                      	#Salva 9 no endereço 2 da RAM (Limite das centenas)
tmp(141) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(142) := x"1" & "00" & '1' & x"61";	-- LDA @353                    	#Carrega o valor do KEY1 no acumulador
tmp(143) := x"8" & "00" & '0' & x"3E";	-- CEQ @62                     	#Compara o valor do KEY1 com 62 (0)
tmp(144) := x"7" & "00" & '0' & x"78";	-- JEQ @120           	#Se o valor do KEY1 for 0 (nao setou o limite das centenas), vai para o label LimCen (Limite das centenas)
tmp(145) := x"5" & "00" & '1' & x"FE";	-- STA @510                    	#Limpa leitura KEY1
tmp(146) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(147) := x"1" & "00" & '1' & x"40";	-- LDA @320                    	#Carrega valor das chaves SW0 a SW7 no acumulador
tmp(148) := x"8" & "00" & '0' & x"14";	-- CEQ @20                     	#Compara o valor das chaves SW0 a SW7 com 20 (10)
tmp(149) := x"7" & "00" & '0' & x"A3";	-- JEQ @163           	#Se o valor das chaves SW0 a SW7 for 10, vai para o label maxMil (Limite maximo dos milhares)
tmp(150) := x"8" & "00" & '0' & x"15";	-- CEQ @21                     	#Compara o valor das chaves SW0 a SW7 com 21 (11)
tmp(151) := x"7" & "00" & '0' & x"A3";	-- JEQ @163           	#Se o valor das chaves SW0 a SW7 for 11, vai para o label maxMil (Limite maximo dos milhares)
tmp(152) := x"8" & "00" & '0' & x"16";	-- CEQ @22                     	#Compara o valor das chaves SW0 a SW7 com 22 (12)
tmp(153) := x"7" & "00" & '0' & x"A3";	-- JEQ @163           	#Se o valor das chaves SW0 a SW7 for 12, vai para o label maxMil (Limite maximo dos milhares)
tmp(154) := x"8" & "00" & '0' & x"17";	-- CEQ @23                     	#Compara o valor das chaves SW0 a SW7 com 23 (13)
tmp(155) := x"7" & "00" & '0' & x"A3";	-- JEQ @163           	#Se o valor das chaves SW0 a SW7 for 13, vai para o label maxMil (Limite maximo dos milhares)
tmp(156) := x"8" & "00" & '0' & x"18";	-- CEQ @24                     	#Compara o valor das chaves SW0 a SW7 com 24 (14)
tmp(157) := x"7" & "00" & '0' & x"A3";	-- JEQ @163           	#Se o valor das chaves SW0 a SW7 for 14, vai para o label maxMil (Limite maximo dos milhares)
tmp(158) := x"8" & "00" & '0' & x"19";	-- CEQ @25                     	#Compara o valor das chaves SW0 a SW7 com 25 (15)
tmp(159) := x"7" & "00" & '0' & x"A3";	-- JEQ @163           	#Se o valor das chaves SW0 a SW7 for 15, vai para o label maxMil (Limite maximo dos milhares)
tmp(160) := x"5" & "00" & '1' & x"23";	-- STA @291                    	#Mostra o valor do acumulador HEX 3 (milhares)
tmp(161) := x"5" & "00" & '0' & x"03";	-- STA @3                      	#Salva o valor do acumulador no endereço 3 da RAM (Limite dos milhares)
tmp(162) := x"6" & "00" & '0' & x"A7";	-- JMP @167           	#Vai para o label MILOK (Milhares menor que o limite)
tmp(163) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(164) := x"1" & "00" & '0' & x"13";	-- LDA @19                     	#Carrega 19 no acumulador
tmp(165) := x"5" & "00" & '1' & x"23";	-- STA @291                    	#Mostra o valor do acumulador HEX 3 (milhares)
tmp(166) := x"5" & "00" & '0' & x"03";	-- STA @3                      	#Salva 9 no endereço 3 da RAM (Limite dos milhares)
tmp(167) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(168) := x"1" & "00" & '1' & x"61";	-- LDA @353                    	#Carrega o valor do KEY1 no acumulador
tmp(169) := x"8" & "00" & '0' & x"3E";	-- CEQ @62                     	#Compara o valor do KEY1 com 62 (0)
tmp(170) := x"7" & "00" & '0' & x"92";	-- JEQ @146           	#Se o valor do KEY1 for 0 (nao setou o limite dos milhares), vai para o label LimMil (Limite dos milhares)
tmp(171) := x"5" & "00" & '1' & x"FE";	-- STA @510                    	#Limpa leitura KEY1
tmp(172) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(173) := x"1" & "00" & '1' & x"40";	-- LDA @320                    	#Carrega valor das chaves SW0 a SW7 no acumulador
tmp(174) := x"8" & "00" & '0' & x"14";	-- CEQ @20                     	#Compara o valor das chaves SW0 a SW7 com 20 (10)
tmp(175) := x"7" & "00" & '0' & x"BD";	-- JEQ @189           	#Se o valor das chaves SW0 a SW7 for 10, vai para o label maxDezM (Limite maximo das dezenas de milhares)
tmp(176) := x"8" & "00" & '0' & x"15";	-- CEQ @21                     	#Compara o valor das chaves SW0 a SW7 com 21 (11)
tmp(177) := x"7" & "00" & '0' & x"BD";	-- JEQ @189           	#Se o valor das chaves SW0 a SW7 for 11, vai para o label maxDezM (Limite maximo das dezenas de milhares)
tmp(178) := x"8" & "00" & '0' & x"16";	-- CEQ @22                     	#Compara o valor das chaves SW0 a SW7 com 22 (12)
tmp(179) := x"7" & "00" & '0' & x"BD";	-- JEQ @189           	#Se o valor das chaves SW0 a SW7 for 12, vai para o label maxDezM (Limite maximo das dezenas de milhares)
tmp(180) := x"8" & "00" & '0' & x"17";	-- CEQ @23                     	#Compara o valor das chaves SW0 a SW7 com 23 (13)
tmp(181) := x"7" & "00" & '0' & x"BD";	-- JEQ @189           	#Se o valor das chaves SW0 a SW7 for 13, vai para o label maxDezM (Limite maximo das dezenas de milhares)
tmp(182) := x"8" & "00" & '0' & x"18";	-- CEQ @24                     	#Compara o valor das chaves SW0 a SW7 com 24 (14)
tmp(183) := x"7" & "00" & '0' & x"BD";	-- JEQ @189           	#Se o valor das chaves SW0 a SW7 for 14, vai para o label maxDezM (Limite maximo das dezenas de milhares)
tmp(184) := x"8" & "00" & '0' & x"19";	-- CEQ @25                     	#Compara o valor das chaves SW0 a SW7 com 25 (15)
tmp(185) := x"7" & "00" & '0' & x"BD";	-- JEQ @189           	#Se o valor das chaves SW0 a SW7 for 15, vai para o label maxDezM (Limite maximo das dezenas de milhares)
tmp(186) := x"5" & "00" & '1' & x"24";	-- STA @292                    	#Mostra o valor do acumulador HEX 4 (dezenas de milhares)
tmp(187) := x"5" & "00" & '0' & x"04";	-- STA @4                      	#Salva o valor do acumulador no endereço 4 da RAM (Limite das dezenas de milhares)
tmp(188) := x"6" & "00" & '0' & x"C1";	-- JMP @193           	#Vai para o label DEZMOK (Dezenas de milhares menor que o limite)
tmp(189) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(190) := x"1" & "00" & '0' & x"13";	-- LDA @19                     	#Carrega 19 no acumulador
tmp(191) := x"5" & "00" & '1' & x"24";	-- STA @292                    	#Mostra o valor do acumulador HEX 4 (dezenas de milhares)
tmp(192) := x"5" & "00" & '0' & x"04";	-- STA @4                      	#Salva 9 no endereço 4 da RAM (Limite das dezenas de milhares)
tmp(193) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(194) := x"1" & "00" & '1' & x"61";	-- LDA @353                    	#Carrega o valor do KEY1 no acumulador
tmp(195) := x"8" & "00" & '0' & x"3E";	-- CEQ @62                     	#Compara o valor do KEY1 com 62 (0)
tmp(196) := x"7" & "00" & '0' & x"AC";	-- JEQ @172           	#Se o valor do KEY1 for 0 (nao setou o limite das dezenas de milhares), vai para o label LimDezM (Limite das dezenas de milhares)
tmp(197) := x"5" & "00" & '1' & x"FE";	-- STA @510                    	#Limpa leitura KEY1
tmp(198) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(199) := x"1" & "00" & '1' & x"40";	-- LDA @320                    	#Carrega valor das chaves SW0 a SW7 no acumulador
tmp(200) := x"8" & "00" & '0' & x"14";	-- CEQ @20                     	#Compara o valor das chaves SW0 a SW7 com 20 (10)
tmp(201) := x"7" & "00" & '0' & x"D7";	-- JEQ @215           	#Se o valor das chaves SW0 a SW7 for 10, vai para o label maxCenM (Limite maximo das centenas de milhares)
tmp(202) := x"8" & "00" & '0' & x"15";	-- CEQ @21                     	#Compara o valor das chaves SW0 a SW7 com 21 (11)
tmp(203) := x"7" & "00" & '0' & x"D7";	-- JEQ @215           	#Se o valor das chaves SW0 a SW7 for 11, vai para o label maxCenM (Limite maximo das centenas de milhares)
tmp(204) := x"8" & "00" & '0' & x"16";	-- CEQ @22                     	#Compara o valor das chaves SW0 a SW7 com 22 (12)
tmp(205) := x"7" & "00" & '0' & x"D7";	-- JEQ @215           	#Se o valor das chaves SW0 a SW7 for 12, vai para o label maxCenM (Limite maximo das centenas de milhares)
tmp(206) := x"8" & "00" & '0' & x"17";	-- CEQ @23                     	#Compara o valor das chaves SW0 a SW7 com 23 (13)
tmp(207) := x"7" & "00" & '0' & x"D7";	-- JEQ @215           	#Se o valor das chaves SW0 a SW7 for 13, vai para o label maxCenM (Limite maximo das centenas de milhares)
tmp(208) := x"8" & "00" & '0' & x"18";	-- CEQ @24                     	#Compara o valor das chaves SW0 a SW7 com 24 (14)
tmp(209) := x"7" & "00" & '0' & x"D7";	-- JEQ @215           	#Se o valor das chaves SW0 a SW7 for 14, vai para o label maxCenM (Limite maximo das centenas de milhares)
tmp(210) := x"8" & "00" & '0' & x"19";	-- CEQ @25                     	#Compara o valor das chaves SW0 a SW7 com 25 (15)
tmp(211) := x"7" & "00" & '0' & x"D7";	-- JEQ @215           	#Se o valor das chaves SW0 a SW7 for 15, vai para o label maxCenM (Limite maximo das centenas de milhares)
tmp(212) := x"5" & "00" & '1' & x"25";	-- STA @293                    	#Mostra o valor do acumulador HEX 5 (centenas de milhares)
tmp(213) := x"5" & "00" & '0' & x"05";	-- STA @5                      	#Salva o valor do acumulador no endereço 5 da RAM (Limite das centenas de milhares)
tmp(214) := x"6" & "00" & '0' & x"DB";	-- JMP @219           	#Vai para o label CENMOK (Centenas de milhares menor que o limite)
tmp(215) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(216) := x"1" & "00" & '0' & x"13";	-- LDA @19                     	#Carrega 19 no acumulador
tmp(217) := x"5" & "00" & '1' & x"25";	-- STA @293                    	#Mostra o valor do acumulador HEX 5 (centenas de milhares)
tmp(218) := x"5" & "00" & '0' & x"05";	-- STA @5                      	#Salva 9 no endereço 5 da RAM (Limite das centenas de milhares)
tmp(219) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(220) := x"1" & "00" & '1' & x"61";	-- LDA @353                    	#Carrega o valor do KEY1 no acumulador
tmp(221) := x"8" & "00" & '0' & x"3E";	-- CEQ @62                     	#Compara o valor do KEY1 com 62 (0)
tmp(222) := x"7" & "00" & '0' & x"C6";	-- JEQ @198           	#Se o valor do KEY1 for 0 (nao setou o limite das centenas de milhares), vai para o label LimCenM (Limite das centenas de milhares)
tmp(223) := x"5" & "00" & '1' & x"FE";	-- STA @510                    	#Limpa leitura KEY1
tmp(224) := x"1" & "00" & '0' & x"0A";	-- LDA @10                     	#Carrega o valor do endereço 10 da RAM no acumulador (valor atual das unidades)
tmp(225) := x"5" & "00" & '1' & x"20";	-- STA @288                    	#Mostra o valor do acumulador HEX 0 (unidades)
tmp(226) := x"1" & "00" & '0' & x"0B";	-- LDA @11                     	#Carrega o valor do endereço 11 da RAM no acumulador (valor atual das dezenas)
tmp(227) := x"5" & "00" & '1' & x"21";	-- STA @289                    	#Mostra o valor do acumulador HEX 1 (dezenas)
tmp(228) := x"1" & "00" & '0' & x"0C";	-- LDA @12                     	#Carrega o valor do endereço 12 da RAM no acumulador (valor atual das centenas)
tmp(229) := x"5" & "00" & '1' & x"22";	-- STA @290                    	#Mostra o valor do acumulador HEX 2 (centenas)
tmp(230) := x"1" & "00" & '0' & x"0D";	-- LDA @13                     	#Carrega o valor do endereço 13 da RAM no acumulador (valor atual dos milhares)
tmp(231) := x"5" & "00" & '1' & x"23";	-- STA @291                    	#Mostra o valor do acumulador HEX 3 (milhares)
tmp(232) := x"1" & "00" & '0' & x"0E";	-- LDA @14                     	#Carrega o valor do endereço 14 da RAM no acumulador (valor atual das dezenas de milhares)
tmp(233) := x"5" & "00" & '1' & x"24";	-- STA @292                    	#Mostra o valor do acumulador HEX 4 (dezenas de milhares)
tmp(234) := x"1" & "00" & '0' & x"0F";	-- LDA @15                     	#Carrega o valor do endereço 15 da RAM no acumulador (valor atual das centenas de milhares)
tmp(235) := x"5" & "00" & '1' & x"25";	-- STA @293                    	#Mostra o valor do acumulador HEX 5 (centenas de milhares)
tmp(236) := x"6" & "00" & '0' & x"2B";	-- JMP @43           	#Volta para o label Start (inicio do programa)
tmp(237) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(238) := x"5" & "00" & '1' & x"FF";	-- STA @511                    	#Limpa leitura KEY0
tmp(239) := x"1" & "00" & '0' & x"0A";	-- LDA @10                     	#Carrega o valor do endereço 10 da RAM no acumulador (valor atual das unidades)
tmp(240) := x"2" & "00" & '0' & x"3F";	-- SOMA @63                    	#Soma o valor do acumulador com 63 (1)
tmp(241) := x"8" & "00" & '0' & x"14";	-- CEQ @20                     	#Compara o valor do acumulador com o endereco 20 da RAM (10)
tmp(242) := x"7" & "00" & '0' & x"F5";	-- JEQ @245           	#Se o valor do acumulador for 10, vai para o label IncDez (Incremento das dezenas)
tmp(243) := x"5" & "00" & '0' & x"0A";	-- STA @10                     	#Se o valor do acumulador nao for 10, salva o valor do acumulador no endereço 10 da RAM (valor atual das unidades)
tmp(244) := x"6" & "00" & '1' & x"22";	-- JMP @290           	#Vai para o label Display (Mostra o valor atual)
tmp(245) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(246) := x"1" & "00" & '0' & x"3E";	-- LDA @62                     	#Carrega o valor 62 (0) no acumulador
tmp(247) := x"5" & "00" & '0' & x"0A";	-- STA @10                     	#Zera o valor atual das unidades
tmp(248) := x"1" & "00" & '0' & x"0B";	-- LDA @11                     	#Carrega o valor do endereço 11 da RAM no acumulador (valor atual das dezenas)
tmp(249) := x"2" & "00" & '0' & x"3F";	-- SOMA @63                    	#Soma o valor do acumulador com 63 (1)
tmp(250) := x"8" & "00" & '0' & x"14";	-- CEQ @20                     	#Compara o valor do acumulador com o endereco 20 da RAM (10)
tmp(251) := x"7" & "00" & '0' & x"FE";	-- JEQ @254           	#Se o valor do acumulador for 10, vai para o label IncCen (Incremento das centenas)
tmp(252) := x"5" & "00" & '0' & x"0B";	-- STA @11                     	#Se o valor do acumulador nao for 10, salva o valor do acumulador no endereço 11 da RAM (valor atual das dezenas)
tmp(253) := x"6" & "00" & '1' & x"22";	-- JMP @290           	#Vai para o label Display (Mostra o valor atual)
tmp(254) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(255) := x"1" & "00" & '0' & x"3E";	-- LDA @62                     	#Carrega o valor 62 (0) no acumulador
tmp(256) := x"5" & "00" & '0' & x"0B";	-- STA @11                     	#Zera o valor atual das dezenas
tmp(257) := x"1" & "00" & '0' & x"0C";	-- LDA @12                     	#Carrega o valor do endereço 12 da RAM no acumulador (valor atual das centenas)
tmp(258) := x"2" & "00" & '0' & x"3F";	-- SOMA @63                    	#Soma o valor do acumulador com 63 (1)
tmp(259) := x"8" & "00" & '0' & x"14";	-- CEQ @20                     	#Compara o valor do acumulador com o endereco 20 da RAM (10)
tmp(260) := x"7" & "00" & '1' & x"07";	-- JEQ @263           	#Se o valor do acumulador for 10, vai para o label IncMil (Incremento dos milhares)
tmp(261) := x"5" & "00" & '0' & x"0C";	-- STA @12                     	#Se o valor do acumulador nao for 10, salva o valor do acumulador no endereço 12 da RAM (valor atual das centenas)
tmp(262) := x"6" & "00" & '1' & x"22";	-- JMP @290           	#Vai para o label Display (Mostra o valor atual)
tmp(263) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(264) := x"1" & "00" & '0' & x"3E";	-- LDA @62                     	#Carrega o valor 62 (0) no acumulador
tmp(265) := x"5" & "00" & '0' & x"0C";	-- STA @12                     	#Zera o valor atual das centenas
tmp(266) := x"1" & "00" & '0' & x"0D";	-- LDA @13                     	#Carrega o valor do endereço 13 da RAM no acumulador (valor atual dos milhares)
tmp(267) := x"2" & "00" & '0' & x"3F";	-- SOMA @63                    	#Soma o valor do acumulador com 63 (1)
tmp(268) := x"8" & "00" & '0' & x"14";	-- CEQ @20                     	#Compara o valor do acumulador com o endereco 20 da RAM (10)
tmp(269) := x"7" & "00" & '1' & x"10";	-- JEQ @272           	#Se o valor do acumulador for 10, vai para o label IncDezM (Incremento das dezenas de milhares)
tmp(270) := x"5" & "00" & '0' & x"0D";	-- STA @13                     	#Se o valor do acumulador nao for 10, salva o valor do acumulador no endereço 13 da RAM (valor atual dos milhares)
tmp(271) := x"6" & "00" & '1' & x"22";	-- JMP @290           	#Vai para o label Display (Mostra o valor atual)
tmp(272) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(273) := x"1" & "00" & '0' & x"3E";	-- LDA @62                     	#Carrega o valor 62 (0) no acumulador
tmp(274) := x"5" & "00" & '0' & x"0D";	-- STA @13                     	#Zera o valor atual dos milhares
tmp(275) := x"1" & "00" & '0' & x"0E";	-- LDA @14                     	#Carrega o valor do endereço 14 da RAM no acumulador (valor atual das dezenas de milhares)
tmp(276) := x"2" & "00" & '0' & x"3F";	-- SOMA @63                    	#Soma o valor do acumulador com 63 (1)
tmp(277) := x"8" & "00" & '0' & x"14";	-- CEQ @20                     	#Compara o valor do acumulador com o endereco 20 da RAM (10)
tmp(278) := x"7" & "00" & '1' & x"19";	-- JEQ @281           	#Se o valor do acumulador for 10, vai para o label IncCenM (Incremento das centenas de milhares)
tmp(279) := x"5" & "00" & '0' & x"0E";	-- STA @14                     	#Se o valor do acumulador nao for 10, salva o valor do acumulador no endereço 14 da RAM (valor atual das dezenas de milhares)
tmp(280) := x"6" & "00" & '1' & x"22";	-- JMP @290           	#Vai para o label Display (Mostra o valor atual)
tmp(281) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(282) := x"1" & "00" & '0' & x"3E";	-- LDA @62                     	#Carrega o valor 62 (0) no acumulador
tmp(283) := x"5" & "00" & '0' & x"0E";	-- STA @14                     	#Zera o valor atual das dezenas de milhares
tmp(284) := x"1" & "00" & '0' & x"0F";	-- LDA @15                     	#Carrega o valor do endereço 15 da RAM no acumulador (valor atual das centenas de milhares)
tmp(285) := x"2" & "00" & '0' & x"3F";	-- SOMA @63                    	#Soma o valor do acumulador com 63 (1)
tmp(286) := x"8" & "00" & '0' & x"14";	-- CEQ @20                     	#Compara o valor do acumulador com o endereco 20 da RAM (10)
tmp(287) := x"7" & "00" & '1' & x"30";	-- JEQ @304           	#Se o valor do acumulador for 10, vai para o label NoveNove (valor nos displays igual a 999999)
tmp(288) := x"5" & "00" & '0' & x"0F";	-- STA @15                     	#Se o valor do acumulador nao for 10, salva o valor do acumulador no endereço 15 da RAM (valor atual das centenas de milhares)
tmp(289) := x"6" & "00" & '1' & x"22";	-- JMP @290           	#Vai para o label Display (Mostra o valor atual)
tmp(290) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(291) := x"1" & "00" & '0' & x"0A";	-- LDA @10                     	#Carrega o valor do endereço 10 da RAM no acumulador (valor atual das unidades)
tmp(292) := x"5" & "00" & '1' & x"20";	-- STA @288                    	#Salva o valor do acumulador no HEX 0
tmp(293) := x"1" & "00" & '0' & x"0B";	-- LDA @11                     	#Carrega o valor do endereço 11 da RAM no acumulador (valor atual das dezenas)
tmp(294) := x"5" & "00" & '1' & x"21";	-- STA @289                    	#Salva o valor do acumulador no HEX 1
tmp(295) := x"1" & "00" & '0' & x"0C";	-- LDA @12                     	#Carrega o valor do endereço 12 da RAM no acumulador (valor atual das centenas)
tmp(296) := x"5" & "00" & '1' & x"22";	-- STA @290                    	#Salva o valor do acumulador no HEX 2
tmp(297) := x"1" & "00" & '0' & x"0D";	-- LDA @13                     	#Carrega o valor do endereço 13 da RAM no acumulador (valor atual dos milhares)
tmp(298) := x"5" & "00" & '1' & x"23";	-- STA @291                    	#Salva o valor do acumulador no HEX 3
tmp(299) := x"1" & "00" & '0' & x"0E";	-- LDA @14                     	#Carrega o valor do endereço 14 da RAM no acumulador (valor atual das dezenas de milhares)
tmp(300) := x"5" & "00" & '1' & x"24";	-- STA @292                    	#Salva o valor do acumulador no HEX 4
tmp(301) := x"1" & "00" & '0' & x"0F";	-- LDA @15                     	#Carrega o valor do endereço 15 da RAM no acumulador (valor atual das centenas de milhares)
tmp(302) := x"5" & "00" & '1' & x"25";	-- STA @293                    	#Salva o valor do acumulador no HEX 5
tmp(303) := x"6" & "00" & '1' & x"37";	-- JMP @311           	#Vai para o label CompLim (Compara o valor atual com o valor do limite)
tmp(304) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(305) := x"1" & "00" & '0' & x"3F";	-- LDA @63                     	#Carrega o valor 63 (1) no acumulador
tmp(306) := x"5" & "00" & '1' & x"02";	-- STA @258                    	#Ascende o LED 9
tmp(307) := x"1" & "00" & '1' & x"64";	-- LDA @356                    	#Carrega o valor do Reset no acumulador
tmp(308) := x"8" & "00" & '0' & x"3F";	-- CEQ @63                     	#Compara o valor do acumulador com 63 (1)
tmp(309) := x"7" & "00" & '0' & x"00";	-- JEQ @0           	#Se o valor do acumulador for 1, vai para o label Reset (Reseta o programa)
tmp(310) := x"6" & "00" & '1' & x"30";	-- JMP @304           	#Se o valor do acumulador nao for 1, vai para o label NoveNove
tmp(311) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(312) := x"1" & "00" & '0' & x"0A";	-- LDA @10                     	#Carrega o valor do endereço 10 da RAM no acumulador (valor atual das unidades)
tmp(313) := x"8" & "00" & '0' & x"00";	-- CEQ @0                      	#Compara o valor do acumulador com o endereco 0 da RAM (limite das unidades)
tmp(314) := x"7" & "00" & '1' & x"3C";	-- JEQ @316           	#Se for igual, vai para o label CompDez (Compara o valor atual das dezenas com o valor do limite das dezenas)
tmp(315) := x"6" & "00" & '0' & x"2B";	-- JMP @43           	#Se nao for igual, vai para o label Start (Loop principal)
tmp(316) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(317) := x"1" & "00" & '0' & x"0B";	-- LDA @11                     	#Carrega o valor do endereço 11 da RAM no acumulador (valor atual das dezenas)
tmp(318) := x"8" & "00" & '0' & x"01";	-- CEQ @1                      	#Compara o valor do acumulador com o endereco 1 da RAM (limite das dezenas)
tmp(319) := x"7" & "00" & '1' & x"41";	-- JEQ @321           	#Se for igual, vai para o label CompCen (Compara o valor atual das centenas com o valor do limite das centenas)
tmp(320) := x"6" & "00" & '0' & x"2B";	-- JMP @43           	#Se nao for igual, vai para o label Start (Loop principal)
tmp(321) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(322) := x"1" & "00" & '0' & x"0C";	-- LDA @12                     	#Carrega o valor do endereço 12 da RAM no acumulador (valor atual das centenas)
tmp(323) := x"8" & "00" & '0' & x"02";	-- CEQ @2                      	#Compara o valor do acumulador com o endereco 2 da RAM (limite das centenas)
tmp(324) := x"7" & "00" & '1' & x"46";	-- JEQ @326           	#Se for igual, vai para o label CompMil (Compara o valor atual dos milhares com o valor do limite dos milhares)
tmp(325) := x"6" & "00" & '0' & x"2B";	-- JMP @43           	#Se nao for igual, vai para o label Start (Loop principal)
tmp(326) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(327) := x"1" & "00" & '0' & x"0D";	-- LDA @13                     	#Carrega o valor do endereço 13 da RAM no acumulador (valor atual dos milhares)
tmp(328) := x"8" & "00" & '0' & x"03";	-- CEQ @3                      	#Compara o valor do acumulador com o endereco 3 da RAM (limite dos milhares)
tmp(329) := x"7" & "00" & '1' & x"4B";	-- JEQ @331           	#Se for igual, vai para o label CompDezM (Compara o valor atual das dezenas de milhares com o valor do limite das dezenas de milhares)
tmp(330) := x"6" & "00" & '0' & x"2B";	-- JMP @43           	#Se nao for igual, vai para o label Start (Loop principal)
tmp(331) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(332) := x"1" & "00" & '0' & x"0E";	-- LDA @14                     	#Carrega o valor do endereço 14 da RAM no acumulador (valor atual das dezenas de milhares)
tmp(333) := x"8" & "00" & '0' & x"04";	-- CEQ @4                      	#Compara o valor do acumulador com o endereco 4 da RAM (limite das dezenas de milhares)
tmp(334) := x"7" & "00" & '1' & x"50";	-- JEQ @336           	#Se for igual, vai para o label CompCenM (Compara o valor atual das centenas de milhares com o valor do limite das centenas de milhares)
tmp(335) := x"6" & "00" & '0' & x"2B";	-- JMP @43           	#Se nao for igual, vai para o label Start (Loop principal)
tmp(336) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(337) := x"1" & "00" & '0' & x"0F";	-- LDA @15                     	#Carrega o valor do endereço 15 da RAM no acumulador (valor atual das centenas de milhares)
tmp(338) := x"8" & "00" & '0' & x"05";	-- CEQ @5                      	#Compara o valor do acumulador com o endereco 5 da RAM (limite das centenas de milhares)
tmp(339) := x"7" & "00" & '1' & x"55";	-- JEQ @341           	#Se for igual, vai para o label Fim (Fim do programa)
tmp(340) := x"6" & "00" & '0' & x"2B";	-- JMP @43           	#Se nao for igual, vai para o label Start (Loop principal)
tmp(341) := x"0" & "00" & '0' & x"00";	-- NOP
tmp(342) := x"1" & "00" & '0' & x"3F";	-- LDA @63                     	#Carrega o valor 63 (1) no acumulador
tmp(343) := x"5" & "00" & '1' & x"02";	-- STA @258                    	#Ascende o LED 9
tmp(344) := x"5" & "00" & '1' & x"01";	-- STA @257                    	#Ascende o LED 8
tmp(345) := x"4" & "00" & '0' & x"FF";	-- LDI $255                    	#Carrega o valor 255 no acumulador
tmp(346) := x"5" & "00" & '1' & x"00";	-- STA @256                    	#Ascende os LEDs 7 a 0
tmp(347) := x"1" & "00" & '1' & x"64";	-- LDA @356                    	#Carrega o valor do Reset no acumulador
tmp(348) := x"8" & "00" & '0' & x"3F";	-- CEQ @63                     	#Compara o valor do acumulador com 63 (1)
tmp(349) := x"7" & "00" & '0' & x"00";	-- JEQ @0           	#Se o valor do acumulador for 1, vai para o label Reset (Reseta o programa)
tmp(350) := x"6" & "00" & '1' & x"55";	-- JMP @341           	#Se o valor do acumulador nao for 1, vai para o label Fim



        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;